// finalProject.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module finalProject (
		output wire [9:0]  a0_external_connection_export,           //           a0_external_connection.export
		output wire [9:0]  a1_external_connection_export,           //           a1_external_connection.export
		output wire [9:0]  a2_external_connection_export,           //           a2_external_connection.export
		output wire [9:0]  a3_external_connection_export,           //           a3_external_connection.export
		output wire [15:0] amp_export,                              //                              amp.export
		input  wire        clk_clk,                                 //                              clk.clk
		output wire [9:0]  d0_external_connection_export,           //           d0_external_connection.export
		output wire [9:0]  d1_external_connection_export,           //           d1_external_connection.export
		output wire [9:0]  d2_external_connection_export,           //           d2_external_connection.export
		output wire [9:0]  d3_external_connection_export,           //           d3_external_connection.export
		output wire [15:0] hex_digits_export,                       //                       hex_digits.export
		input  wire        i2c_serial_sda_in,                       //                       i2c_serial.sda_in
		input  wire        i2c_serial_scl_in,                       //                                 .scl_in
		output wire        i2c_serial_sda_oe,                       //                                 .sda_oe
		output wire        i2c_serial_scl_oe,                       //                                 .scl_oe
		input  wire [1:0]  key_external_connection_export,          //          key_external_connection.export
		output wire [7:0]  keycode_export,                          //                          keycode.export
		output wire [7:0]  keycode1_export,                         //                         keycode1.export
		output wire [7:0]  keycode2_export,                         //                         keycode2.export
		output wire [7:0]  keycode3_export,                         //                         keycode3.export
		output wire [13:0] leds_export,                             //                             leds.export
		output wire [7:0]  oct_external_connection_export,          //          oct_external_connection.export
		output wire [31:0] phase_incr0_external_connection_export,  //  phase_incr0_external_connection.export
		output wire [31:0] phase_incr10_external_connection_export, // phase_incr10_external_connection.export
		output wire [31:0] phase_incr11_external_connection_export, // phase_incr11_external_connection.export
		output wire [31:0] phase_incr12_external_connection_export, // phase_incr12_external_connection.export
		output wire [31:0] phase_incr13_external_connection_export, // phase_incr13_external_connection.export
		output wire [31:0] phase_incr14_external_connection_export, // phase_incr14_external_connection.export
		output wire [31:0] phase_incr15_external_connection_export, // phase_incr15_external_connection.export
		output wire [31:0] phase_incr16_external_connection_export, // phase_incr16_external_connection.export
		output wire [31:0] phase_incr17_external_connection_export, // phase_incr17_external_connection.export
		output wire [31:0] phase_incr1_external_connection_export,  //  phase_incr1_external_connection.export
		output wire [31:0] phase_incr2_external_connection_export,  //  phase_incr2_external_connection.export
		output wire [31:0] phase_incr3_external_connection_export,  //  phase_incr3_external_connection.export
		output wire [31:0] phase_incr4_external_connection_export,  //  phase_incr4_external_connection.export
		output wire [31:0] phase_incr5_external_connection_export,  //  phase_incr5_external_connection.export
		output wire [31:0] phase_incr6_external_connection_export,  //  phase_incr6_external_connection.export
		output wire [31:0] phase_incr7_external_connection_export,  //  phase_incr7_external_connection.export
		output wire [31:0] phase_incr8_external_connection_export,  //  phase_incr8_external_connection.export
		output wire [31:0] phase_incr9_external_connection_export,  //  phase_incr9_external_connection.export
		output wire [9:0]  r0_external_connection_export,           //           r0_external_connection.export
		output wire [9:0]  r1_external_connection_export,           //           r1_external_connection.export
		output wire [9:0]  r2_external_connection_export,           //           r2_external_connection.export
		output wire [9:0]  r3_external_connection_export,           //           r3_external_connection.export
		input  wire        reset_reset_n,                           //                            reset.reset_n
		output wire [9:0]  s0_external_connection_export,           //           s0_external_connection.export
		output wire [9:0]  s1_external_connection_export,           //           s1_external_connection.export
		output wire [9:0]  s2_external_connection_export,           //           s2_external_connection.export
		output wire [9:0]  s3_external_connection_export,           //           s3_external_connection.export
		output wire        sdram_clk_clk,                           //                        sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                         //                       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                           //                                 .ba
		output wire        sdram_wire_cas_n,                        //                                 .cas_n
		output wire        sdram_wire_cke,                          //                                 .cke
		output wire        sdram_wire_cs_n,                         //                                 .cs_n
		inout  wire [15:0] sdram_wire_dq,                           //                                 .dq
		output wire [1:0]  sdram_wire_dqm,                          //                                 .dqm
		output wire        sdram_wire_ras_n,                        //                                 .ras_n
		output wire        sdram_wire_we_n,                         //                                 .we_n
		input  wire        spi0_MISO,                               //                             spi0.MISO
		output wire        spi0_MOSI,                               //                                 .MOSI
		output wire        spi0_SCLK,                               //                                 .SCLK
		output wire        spi0_SS_n,                               //                                 .SS_n
		input  wire [9:0]  switches_external_connection_export,     //     switches_external_connection.export
		input  wire        usb_gpx_export,                          //                          usb_gpx.export
		input  wire        usb_irq_export,                          //                          usb_irq.export
		output wire        usb_rst_export,                          //                          usb_rst.export
		output wire [7:0]  waveform_external_connection_export      //     waveform_external_connection.export
	);

	wire         sdram_pll_c0_clk;                                           // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;      // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;       // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_i2c_0_csr_readdata;                       // i2c_0:readdata -> mm_interconnect_0:i2c_0_csr_readdata
	wire   [3:0] mm_interconnect_0_i2c_0_csr_address;                        // mm_interconnect_0:i2c_0_csr_address -> i2c_0:addr
	wire         mm_interconnect_0_i2c_0_csr_read;                           // mm_interconnect_0:i2c_0_csr_read -> i2c_0:read
	wire         mm_interconnect_0_i2c_0_csr_write;                          // mm_interconnect_0:i2c_0_csr_write -> i2c_0:write
	wire  [31:0] mm_interconnect_0_i2c_0_csr_writedata;                      // mm_interconnect_0:i2c_0_csr_writedata -> i2c_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;             // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;              // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                 // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;            // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_keycode_s1_chipselect;                    // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                      // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                       // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                         // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                     // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire  [31:0] mm_interconnect_0_usb_irq_s1_readdata;                      // usb_irq:readdata -> mm_interconnect_0:usb_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_irq_s1_address;                       // mm_interconnect_0:usb_irq_s1_address -> usb_irq:address
	wire  [31:0] mm_interconnect_0_usb_gpx_s1_readdata;                      // usb_gpx:readdata -> mm_interconnect_0:usb_gpx_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_gpx_s1_address;                       // mm_interconnect_0:usb_gpx_s1_address -> usb_gpx:address
	wire         mm_interconnect_0_usb_rst_s1_chipselect;                    // mm_interconnect_0:usb_rst_s1_chipselect -> usb_rst:chipselect
	wire  [31:0] mm_interconnect_0_usb_rst_s1_readdata;                      // usb_rst:readdata -> mm_interconnect_0:usb_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_rst_s1_address;                       // mm_interconnect_0:usb_rst_s1_address -> usb_rst:address
	wire         mm_interconnect_0_usb_rst_s1_write;                         // mm_interconnect_0:usb_rst_s1_write -> usb_rst:write_n
	wire  [31:0] mm_interconnect_0_usb_rst_s1_writedata;                     // mm_interconnect_0:usb_rst_s1_writedata -> usb_rst:writedata
	wire         mm_interconnect_0_hex_digits_pio_s1_chipselect;             // mm_interconnect_0:hex_digits_pio_s1_chipselect -> hex_digits_pio:chipselect
	wire  [31:0] mm_interconnect_0_hex_digits_pio_s1_readdata;               // hex_digits_pio:readdata -> mm_interconnect_0:hex_digits_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_digits_pio_s1_address;                // mm_interconnect_0:hex_digits_pio_s1_address -> hex_digits_pio:address
	wire         mm_interconnect_0_hex_digits_pio_s1_write;                  // mm_interconnect_0:hex_digits_pio_s1_write -> hex_digits_pio:write_n
	wire  [31:0] mm_interconnect_0_hex_digits_pio_s1_writedata;              // mm_interconnect_0:hex_digits_pio_s1_writedata -> hex_digits_pio:writedata
	wire         mm_interconnect_0_leds_pio_s1_chipselect;                   // mm_interconnect_0:leds_pio_s1_chipselect -> leds_pio:chipselect
	wire  [31:0] mm_interconnect_0_leds_pio_s1_readdata;                     // leds_pio:readdata -> mm_interconnect_0:leds_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_pio_s1_address;                      // mm_interconnect_0:leds_pio_s1_address -> leds_pio:address
	wire         mm_interconnect_0_leds_pio_s1_write;                        // mm_interconnect_0:leds_pio_s1_write -> leds_pio:write_n
	wire  [31:0] mm_interconnect_0_leds_pio_s1_writedata;                    // mm_interconnect_0:leds_pio_s1_writedata -> leds_pio:writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                          // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                           // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_timer_s1_chipselect;                      // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                        // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_s1_address;                         // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                           // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                       // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_phase_incr0_s1_chipselect;                // mm_interconnect_0:phase_incr0_s1_chipselect -> phase_incr0:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr0_s1_readdata;                  // phase_incr0:readdata -> mm_interconnect_0:phase_incr0_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr0_s1_address;                   // mm_interconnect_0:phase_incr0_s1_address -> phase_incr0:address
	wire         mm_interconnect_0_phase_incr0_s1_write;                     // mm_interconnect_0:phase_incr0_s1_write -> phase_incr0:write_n
	wire  [31:0] mm_interconnect_0_phase_incr0_s1_writedata;                 // mm_interconnect_0:phase_incr0_s1_writedata -> phase_incr0:writedata
	wire         mm_interconnect_0_phase_incr1_s1_chipselect;                // mm_interconnect_0:phase_incr1_s1_chipselect -> phase_incr1:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr1_s1_readdata;                  // phase_incr1:readdata -> mm_interconnect_0:phase_incr1_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr1_s1_address;                   // mm_interconnect_0:phase_incr1_s1_address -> phase_incr1:address
	wire         mm_interconnect_0_phase_incr1_s1_write;                     // mm_interconnect_0:phase_incr1_s1_write -> phase_incr1:write_n
	wire  [31:0] mm_interconnect_0_phase_incr1_s1_writedata;                 // mm_interconnect_0:phase_incr1_s1_writedata -> phase_incr1:writedata
	wire         mm_interconnect_0_phase_incr2_s1_chipselect;                // mm_interconnect_0:phase_incr2_s1_chipselect -> phase_incr2:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr2_s1_readdata;                  // phase_incr2:readdata -> mm_interconnect_0:phase_incr2_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr2_s1_address;                   // mm_interconnect_0:phase_incr2_s1_address -> phase_incr2:address
	wire         mm_interconnect_0_phase_incr2_s1_write;                     // mm_interconnect_0:phase_incr2_s1_write -> phase_incr2:write_n
	wire  [31:0] mm_interconnect_0_phase_incr2_s1_writedata;                 // mm_interconnect_0:phase_incr2_s1_writedata -> phase_incr2:writedata
	wire         mm_interconnect_0_phase_incr3_s1_chipselect;                // mm_interconnect_0:phase_incr3_s1_chipselect -> phase_incr3:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr3_s1_readdata;                  // phase_incr3:readdata -> mm_interconnect_0:phase_incr3_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr3_s1_address;                   // mm_interconnect_0:phase_incr3_s1_address -> phase_incr3:address
	wire         mm_interconnect_0_phase_incr3_s1_write;                     // mm_interconnect_0:phase_incr3_s1_write -> phase_incr3:write_n
	wire  [31:0] mm_interconnect_0_phase_incr3_s1_writedata;                 // mm_interconnect_0:phase_incr3_s1_writedata -> phase_incr3:writedata
	wire         mm_interconnect_0_phase_incr4_s1_chipselect;                // mm_interconnect_0:phase_incr4_s1_chipselect -> phase_incr4:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr4_s1_readdata;                  // phase_incr4:readdata -> mm_interconnect_0:phase_incr4_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr4_s1_address;                   // mm_interconnect_0:phase_incr4_s1_address -> phase_incr4:address
	wire         mm_interconnect_0_phase_incr4_s1_write;                     // mm_interconnect_0:phase_incr4_s1_write -> phase_incr4:write_n
	wire  [31:0] mm_interconnect_0_phase_incr4_s1_writedata;                 // mm_interconnect_0:phase_incr4_s1_writedata -> phase_incr4:writedata
	wire         mm_interconnect_0_phase_incr5_s1_chipselect;                // mm_interconnect_0:phase_incr5_s1_chipselect -> phase_incr5:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr5_s1_readdata;                  // phase_incr5:readdata -> mm_interconnect_0:phase_incr5_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr5_s1_address;                   // mm_interconnect_0:phase_incr5_s1_address -> phase_incr5:address
	wire         mm_interconnect_0_phase_incr5_s1_write;                     // mm_interconnect_0:phase_incr5_s1_write -> phase_incr5:write_n
	wire  [31:0] mm_interconnect_0_phase_incr5_s1_writedata;                 // mm_interconnect_0:phase_incr5_s1_writedata -> phase_incr5:writedata
	wire         mm_interconnect_0_phase_incr6_s1_chipselect;                // mm_interconnect_0:phase_incr6_s1_chipselect -> phase_incr6:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr6_s1_readdata;                  // phase_incr6:readdata -> mm_interconnect_0:phase_incr6_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr6_s1_address;                   // mm_interconnect_0:phase_incr6_s1_address -> phase_incr6:address
	wire         mm_interconnect_0_phase_incr6_s1_write;                     // mm_interconnect_0:phase_incr6_s1_write -> phase_incr6:write_n
	wire  [31:0] mm_interconnect_0_phase_incr6_s1_writedata;                 // mm_interconnect_0:phase_incr6_s1_writedata -> phase_incr6:writedata
	wire         mm_interconnect_0_phase_incr7_s1_chipselect;                // mm_interconnect_0:phase_incr7_s1_chipselect -> phase_incr7:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr7_s1_readdata;                  // phase_incr7:readdata -> mm_interconnect_0:phase_incr7_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr7_s1_address;                   // mm_interconnect_0:phase_incr7_s1_address -> phase_incr7:address
	wire         mm_interconnect_0_phase_incr7_s1_write;                     // mm_interconnect_0:phase_incr7_s1_write -> phase_incr7:write_n
	wire  [31:0] mm_interconnect_0_phase_incr7_s1_writedata;                 // mm_interconnect_0:phase_incr7_s1_writedata -> phase_incr7:writedata
	wire         mm_interconnect_0_phase_incr8_s1_chipselect;                // mm_interconnect_0:phase_incr8_s1_chipselect -> phase_incr8:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr8_s1_readdata;                  // phase_incr8:readdata -> mm_interconnect_0:phase_incr8_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr8_s1_address;                   // mm_interconnect_0:phase_incr8_s1_address -> phase_incr8:address
	wire         mm_interconnect_0_phase_incr8_s1_write;                     // mm_interconnect_0:phase_incr8_s1_write -> phase_incr8:write_n
	wire  [31:0] mm_interconnect_0_phase_incr8_s1_writedata;                 // mm_interconnect_0:phase_incr8_s1_writedata -> phase_incr8:writedata
	wire         mm_interconnect_0_phase_incr9_s1_chipselect;                // mm_interconnect_0:phase_incr9_s1_chipselect -> phase_incr9:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr9_s1_readdata;                  // phase_incr9:readdata -> mm_interconnect_0:phase_incr9_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr9_s1_address;                   // mm_interconnect_0:phase_incr9_s1_address -> phase_incr9:address
	wire         mm_interconnect_0_phase_incr9_s1_write;                     // mm_interconnect_0:phase_incr9_s1_write -> phase_incr9:write_n
	wire  [31:0] mm_interconnect_0_phase_incr9_s1_writedata;                 // mm_interconnect_0:phase_incr9_s1_writedata -> phase_incr9:writedata
	wire         mm_interconnect_0_phase_incr10_s1_chipselect;               // mm_interconnect_0:phase_incr10_s1_chipselect -> phase_incr10:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr10_s1_readdata;                 // phase_incr10:readdata -> mm_interconnect_0:phase_incr10_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr10_s1_address;                  // mm_interconnect_0:phase_incr10_s1_address -> phase_incr10:address
	wire         mm_interconnect_0_phase_incr10_s1_write;                    // mm_interconnect_0:phase_incr10_s1_write -> phase_incr10:write_n
	wire  [31:0] mm_interconnect_0_phase_incr10_s1_writedata;                // mm_interconnect_0:phase_incr10_s1_writedata -> phase_incr10:writedata
	wire         mm_interconnect_0_phase_incr11_s1_chipselect;               // mm_interconnect_0:phase_incr11_s1_chipselect -> phase_incr11:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr11_s1_readdata;                 // phase_incr11:readdata -> mm_interconnect_0:phase_incr11_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr11_s1_address;                  // mm_interconnect_0:phase_incr11_s1_address -> phase_incr11:address
	wire         mm_interconnect_0_phase_incr11_s1_write;                    // mm_interconnect_0:phase_incr11_s1_write -> phase_incr11:write_n
	wire  [31:0] mm_interconnect_0_phase_incr11_s1_writedata;                // mm_interconnect_0:phase_incr11_s1_writedata -> phase_incr11:writedata
	wire         mm_interconnect_0_phase_incr12_s1_chipselect;               // mm_interconnect_0:phase_incr12_s1_chipselect -> phase_incr12:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr12_s1_readdata;                 // phase_incr12:readdata -> mm_interconnect_0:phase_incr12_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr12_s1_address;                  // mm_interconnect_0:phase_incr12_s1_address -> phase_incr12:address
	wire         mm_interconnect_0_phase_incr12_s1_write;                    // mm_interconnect_0:phase_incr12_s1_write -> phase_incr12:write_n
	wire  [31:0] mm_interconnect_0_phase_incr12_s1_writedata;                // mm_interconnect_0:phase_incr12_s1_writedata -> phase_incr12:writedata
	wire         mm_interconnect_0_phase_incr13_s1_chipselect;               // mm_interconnect_0:phase_incr13_s1_chipselect -> phase_incr13:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr13_s1_readdata;                 // phase_incr13:readdata -> mm_interconnect_0:phase_incr13_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr13_s1_address;                  // mm_interconnect_0:phase_incr13_s1_address -> phase_incr13:address
	wire         mm_interconnect_0_phase_incr13_s1_write;                    // mm_interconnect_0:phase_incr13_s1_write -> phase_incr13:write_n
	wire  [31:0] mm_interconnect_0_phase_incr13_s1_writedata;                // mm_interconnect_0:phase_incr13_s1_writedata -> phase_incr13:writedata
	wire         mm_interconnect_0_phase_incr14_s1_chipselect;               // mm_interconnect_0:phase_incr14_s1_chipselect -> phase_incr14:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr14_s1_readdata;                 // phase_incr14:readdata -> mm_interconnect_0:phase_incr14_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr14_s1_address;                  // mm_interconnect_0:phase_incr14_s1_address -> phase_incr14:address
	wire         mm_interconnect_0_phase_incr14_s1_write;                    // mm_interconnect_0:phase_incr14_s1_write -> phase_incr14:write_n
	wire  [31:0] mm_interconnect_0_phase_incr14_s1_writedata;                // mm_interconnect_0:phase_incr14_s1_writedata -> phase_incr14:writedata
	wire         mm_interconnect_0_phase_incr15_s1_chipselect;               // mm_interconnect_0:phase_incr15_s1_chipselect -> phase_incr15:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr15_s1_readdata;                 // phase_incr15:readdata -> mm_interconnect_0:phase_incr15_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr15_s1_address;                  // mm_interconnect_0:phase_incr15_s1_address -> phase_incr15:address
	wire         mm_interconnect_0_phase_incr15_s1_write;                    // mm_interconnect_0:phase_incr15_s1_write -> phase_incr15:write_n
	wire  [31:0] mm_interconnect_0_phase_incr15_s1_writedata;                // mm_interconnect_0:phase_incr15_s1_writedata -> phase_incr15:writedata
	wire         mm_interconnect_0_phase_incr16_s1_chipselect;               // mm_interconnect_0:phase_incr16_s1_chipselect -> phase_incr16:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr16_s1_readdata;                 // phase_incr16:readdata -> mm_interconnect_0:phase_incr16_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr16_s1_address;                  // mm_interconnect_0:phase_incr16_s1_address -> phase_incr16:address
	wire         mm_interconnect_0_phase_incr16_s1_write;                    // mm_interconnect_0:phase_incr16_s1_write -> phase_incr16:write_n
	wire  [31:0] mm_interconnect_0_phase_incr16_s1_writedata;                // mm_interconnect_0:phase_incr16_s1_writedata -> phase_incr16:writedata
	wire         mm_interconnect_0_phase_incr17_s1_chipselect;               // mm_interconnect_0:phase_incr17_s1_chipselect -> phase_incr17:chipselect
	wire  [31:0] mm_interconnect_0_phase_incr17_s1_readdata;                 // phase_incr17:readdata -> mm_interconnect_0:phase_incr17_s1_readdata
	wire   [1:0] mm_interconnect_0_phase_incr17_s1_address;                  // mm_interconnect_0:phase_incr17_s1_address -> phase_incr17:address
	wire         mm_interconnect_0_phase_incr17_s1_write;                    // mm_interconnect_0:phase_incr17_s1_write -> phase_incr17:write_n
	wire  [31:0] mm_interconnect_0_phase_incr17_s1_writedata;                // mm_interconnect_0:phase_incr17_s1_writedata -> phase_incr17:writedata
	wire         mm_interconnect_0_keycode1_s1_chipselect;                   // mm_interconnect_0:keycode1_s1_chipselect -> keycode1:chipselect
	wire  [31:0] mm_interconnect_0_keycode1_s1_readdata;                     // keycode1:readdata -> mm_interconnect_0:keycode1_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode1_s1_address;                      // mm_interconnect_0:keycode1_s1_address -> keycode1:address
	wire         mm_interconnect_0_keycode1_s1_write;                        // mm_interconnect_0:keycode1_s1_write -> keycode1:write_n
	wire  [31:0] mm_interconnect_0_keycode1_s1_writedata;                    // mm_interconnect_0:keycode1_s1_writedata -> keycode1:writedata
	wire         mm_interconnect_0_keycode2_s1_chipselect;                   // mm_interconnect_0:keycode2_s1_chipselect -> keycode2:chipselect
	wire  [31:0] mm_interconnect_0_keycode2_s1_readdata;                     // keycode2:readdata -> mm_interconnect_0:keycode2_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode2_s1_address;                      // mm_interconnect_0:keycode2_s1_address -> keycode2:address
	wire         mm_interconnect_0_keycode2_s1_write;                        // mm_interconnect_0:keycode2_s1_write -> keycode2:write_n
	wire  [31:0] mm_interconnect_0_keycode2_s1_writedata;                    // mm_interconnect_0:keycode2_s1_writedata -> keycode2:writedata
	wire         mm_interconnect_0_keycode3_s1_chipselect;                   // mm_interconnect_0:keycode3_s1_chipselect -> keycode3:chipselect
	wire  [31:0] mm_interconnect_0_keycode3_s1_readdata;                     // keycode3:readdata -> mm_interconnect_0:keycode3_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode3_s1_address;                      // mm_interconnect_0:keycode3_s1_address -> keycode3:address
	wire         mm_interconnect_0_keycode3_s1_write;                        // mm_interconnect_0:keycode3_s1_write -> keycode3:write_n
	wire  [31:0] mm_interconnect_0_keycode3_s1_writedata;                    // mm_interconnect_0:keycode3_s1_writedata -> keycode3:writedata
	wire         mm_interconnect_0_amplitude_s1_chipselect;                  // mm_interconnect_0:amplitude_s1_chipselect -> amplitude:chipselect
	wire  [31:0] mm_interconnect_0_amplitude_s1_readdata;                    // amplitude:readdata -> mm_interconnect_0:amplitude_s1_readdata
	wire   [1:0] mm_interconnect_0_amplitude_s1_address;                     // mm_interconnect_0:amplitude_s1_address -> amplitude:address
	wire         mm_interconnect_0_amplitude_s1_write;                       // mm_interconnect_0:amplitude_s1_write -> amplitude:write_n
	wire  [31:0] mm_interconnect_0_amplitude_s1_writedata;                   // mm_interconnect_0:amplitude_s1_writedata -> amplitude:writedata
	wire         mm_interconnect_0_a0_s1_chipselect;                         // mm_interconnect_0:a0_s1_chipselect -> a0:chipselect
	wire  [31:0] mm_interconnect_0_a0_s1_readdata;                           // a0:readdata -> mm_interconnect_0:a0_s1_readdata
	wire   [1:0] mm_interconnect_0_a0_s1_address;                            // mm_interconnect_0:a0_s1_address -> a0:address
	wire         mm_interconnect_0_a0_s1_write;                              // mm_interconnect_0:a0_s1_write -> a0:write_n
	wire  [31:0] mm_interconnect_0_a0_s1_writedata;                          // mm_interconnect_0:a0_s1_writedata -> a0:writedata
	wire         mm_interconnect_0_d0_s1_chipselect;                         // mm_interconnect_0:d0_s1_chipselect -> d0:chipselect
	wire  [31:0] mm_interconnect_0_d0_s1_readdata;                           // d0:readdata -> mm_interconnect_0:d0_s1_readdata
	wire   [1:0] mm_interconnect_0_d0_s1_address;                            // mm_interconnect_0:d0_s1_address -> d0:address
	wire         mm_interconnect_0_d0_s1_write;                              // mm_interconnect_0:d0_s1_write -> d0:write_n
	wire  [31:0] mm_interconnect_0_d0_s1_writedata;                          // mm_interconnect_0:d0_s1_writedata -> d0:writedata
	wire         mm_interconnect_0_s0_s1_chipselect;                         // mm_interconnect_0:s0_s1_chipselect -> s0:chipselect
	wire  [31:0] mm_interconnect_0_s0_s1_readdata;                           // s0:readdata -> mm_interconnect_0:s0_s1_readdata
	wire   [1:0] mm_interconnect_0_s0_s1_address;                            // mm_interconnect_0:s0_s1_address -> s0:address
	wire         mm_interconnect_0_s0_s1_write;                              // mm_interconnect_0:s0_s1_write -> s0:write_n
	wire  [31:0] mm_interconnect_0_s0_s1_writedata;                          // mm_interconnect_0:s0_s1_writedata -> s0:writedata
	wire         mm_interconnect_0_r0_s1_chipselect;                         // mm_interconnect_0:r0_s1_chipselect -> r0:chipselect
	wire  [31:0] mm_interconnect_0_r0_s1_readdata;                           // r0:readdata -> mm_interconnect_0:r0_s1_readdata
	wire   [1:0] mm_interconnect_0_r0_s1_address;                            // mm_interconnect_0:r0_s1_address -> r0:address
	wire         mm_interconnect_0_r0_s1_write;                              // mm_interconnect_0:r0_s1_write -> r0:write_n
	wire  [31:0] mm_interconnect_0_r0_s1_writedata;                          // mm_interconnect_0:r0_s1_writedata -> r0:writedata
	wire         mm_interconnect_0_a1_s1_chipselect;                         // mm_interconnect_0:a1_s1_chipselect -> a1:chipselect
	wire  [31:0] mm_interconnect_0_a1_s1_readdata;                           // a1:readdata -> mm_interconnect_0:a1_s1_readdata
	wire   [1:0] mm_interconnect_0_a1_s1_address;                            // mm_interconnect_0:a1_s1_address -> a1:address
	wire         mm_interconnect_0_a1_s1_write;                              // mm_interconnect_0:a1_s1_write -> a1:write_n
	wire  [31:0] mm_interconnect_0_a1_s1_writedata;                          // mm_interconnect_0:a1_s1_writedata -> a1:writedata
	wire         mm_interconnect_0_d1_s1_chipselect;                         // mm_interconnect_0:d1_s1_chipselect -> d1:chipselect
	wire  [31:0] mm_interconnect_0_d1_s1_readdata;                           // d1:readdata -> mm_interconnect_0:d1_s1_readdata
	wire   [1:0] mm_interconnect_0_d1_s1_address;                            // mm_interconnect_0:d1_s1_address -> d1:address
	wire         mm_interconnect_0_d1_s1_write;                              // mm_interconnect_0:d1_s1_write -> d1:write_n
	wire  [31:0] mm_interconnect_0_d1_s1_writedata;                          // mm_interconnect_0:d1_s1_writedata -> d1:writedata
	wire         mm_interconnect_0_s1_s1_chipselect;                         // mm_interconnect_0:s1_s1_chipselect -> s1:chipselect
	wire  [31:0] mm_interconnect_0_s1_s1_readdata;                           // s1:readdata -> mm_interconnect_0:s1_s1_readdata
	wire   [1:0] mm_interconnect_0_s1_s1_address;                            // mm_interconnect_0:s1_s1_address -> s1:address
	wire         mm_interconnect_0_s1_s1_write;                              // mm_interconnect_0:s1_s1_write -> s1:write_n
	wire  [31:0] mm_interconnect_0_s1_s1_writedata;                          // mm_interconnect_0:s1_s1_writedata -> s1:writedata
	wire         mm_interconnect_0_r1_s1_chipselect;                         // mm_interconnect_0:r1_s1_chipselect -> r1:chipselect
	wire  [31:0] mm_interconnect_0_r1_s1_readdata;                           // r1:readdata -> mm_interconnect_0:r1_s1_readdata
	wire   [1:0] mm_interconnect_0_r1_s1_address;                            // mm_interconnect_0:r1_s1_address -> r1:address
	wire         mm_interconnect_0_r1_s1_write;                              // mm_interconnect_0:r1_s1_write -> r1:write_n
	wire  [31:0] mm_interconnect_0_r1_s1_writedata;                          // mm_interconnect_0:r1_s1_writedata -> r1:writedata
	wire         mm_interconnect_0_a2_s1_chipselect;                         // mm_interconnect_0:a2_s1_chipselect -> a2:chipselect
	wire  [31:0] mm_interconnect_0_a2_s1_readdata;                           // a2:readdata -> mm_interconnect_0:a2_s1_readdata
	wire   [1:0] mm_interconnect_0_a2_s1_address;                            // mm_interconnect_0:a2_s1_address -> a2:address
	wire         mm_interconnect_0_a2_s1_write;                              // mm_interconnect_0:a2_s1_write -> a2:write_n
	wire  [31:0] mm_interconnect_0_a2_s1_writedata;                          // mm_interconnect_0:a2_s1_writedata -> a2:writedata
	wire         mm_interconnect_0_d2_s1_chipselect;                         // mm_interconnect_0:d2_s1_chipselect -> d2:chipselect
	wire  [31:0] mm_interconnect_0_d2_s1_readdata;                           // d2:readdata -> mm_interconnect_0:d2_s1_readdata
	wire   [1:0] mm_interconnect_0_d2_s1_address;                            // mm_interconnect_0:d2_s1_address -> d2:address
	wire         mm_interconnect_0_d2_s1_write;                              // mm_interconnect_0:d2_s1_write -> d2:write_n
	wire  [31:0] mm_interconnect_0_d2_s1_writedata;                          // mm_interconnect_0:d2_s1_writedata -> d2:writedata
	wire         mm_interconnect_0_s2_s1_chipselect;                         // mm_interconnect_0:s2_s1_chipselect -> s2:chipselect
	wire  [31:0] mm_interconnect_0_s2_s1_readdata;                           // s2:readdata -> mm_interconnect_0:s2_s1_readdata
	wire   [1:0] mm_interconnect_0_s2_s1_address;                            // mm_interconnect_0:s2_s1_address -> s2:address
	wire         mm_interconnect_0_s2_s1_write;                              // mm_interconnect_0:s2_s1_write -> s2:write_n
	wire  [31:0] mm_interconnect_0_s2_s1_writedata;                          // mm_interconnect_0:s2_s1_writedata -> s2:writedata
	wire         mm_interconnect_0_r2_s1_chipselect;                         // mm_interconnect_0:r2_s1_chipselect -> r2:chipselect
	wire  [31:0] mm_interconnect_0_r2_s1_readdata;                           // r2:readdata -> mm_interconnect_0:r2_s1_readdata
	wire   [1:0] mm_interconnect_0_r2_s1_address;                            // mm_interconnect_0:r2_s1_address -> r2:address
	wire         mm_interconnect_0_r2_s1_write;                              // mm_interconnect_0:r2_s1_write -> r2:write_n
	wire  [31:0] mm_interconnect_0_r2_s1_writedata;                          // mm_interconnect_0:r2_s1_writedata -> r2:writedata
	wire         mm_interconnect_0_a3_s1_chipselect;                         // mm_interconnect_0:a3_s1_chipselect -> a3:chipselect
	wire  [31:0] mm_interconnect_0_a3_s1_readdata;                           // a3:readdata -> mm_interconnect_0:a3_s1_readdata
	wire   [1:0] mm_interconnect_0_a3_s1_address;                            // mm_interconnect_0:a3_s1_address -> a3:address
	wire         mm_interconnect_0_a3_s1_write;                              // mm_interconnect_0:a3_s1_write -> a3:write_n
	wire  [31:0] mm_interconnect_0_a3_s1_writedata;                          // mm_interconnect_0:a3_s1_writedata -> a3:writedata
	wire         mm_interconnect_0_d3_s1_chipselect;                         // mm_interconnect_0:d3_s1_chipselect -> d3:chipselect
	wire  [31:0] mm_interconnect_0_d3_s1_readdata;                           // d3:readdata -> mm_interconnect_0:d3_s1_readdata
	wire   [1:0] mm_interconnect_0_d3_s1_address;                            // mm_interconnect_0:d3_s1_address -> d3:address
	wire         mm_interconnect_0_d3_s1_write;                              // mm_interconnect_0:d3_s1_write -> d3:write_n
	wire  [31:0] mm_interconnect_0_d3_s1_writedata;                          // mm_interconnect_0:d3_s1_writedata -> d3:writedata
	wire         mm_interconnect_0_s3_s1_chipselect;                         // mm_interconnect_0:s3_s1_chipselect -> s3:chipselect
	wire  [31:0] mm_interconnect_0_s3_s1_readdata;                           // s3:readdata -> mm_interconnect_0:s3_s1_readdata
	wire   [1:0] mm_interconnect_0_s3_s1_address;                            // mm_interconnect_0:s3_s1_address -> s3:address
	wire         mm_interconnect_0_s3_s1_write;                              // mm_interconnect_0:s3_s1_write -> s3:write_n
	wire  [31:0] mm_interconnect_0_s3_s1_writedata;                          // mm_interconnect_0:s3_s1_writedata -> s3:writedata
	wire         mm_interconnect_0_r3_s1_chipselect;                         // mm_interconnect_0:r3_s1_chipselect -> r3:chipselect
	wire  [31:0] mm_interconnect_0_r3_s1_readdata;                           // r3:readdata -> mm_interconnect_0:r3_s1_readdata
	wire   [1:0] mm_interconnect_0_r3_s1_address;                            // mm_interconnect_0:r3_s1_address -> r3:address
	wire         mm_interconnect_0_r3_s1_write;                              // mm_interconnect_0:r3_s1_write -> r3:write_n
	wire  [31:0] mm_interconnect_0_r3_s1_writedata;                          // mm_interconnect_0:r3_s1_writedata -> r3:writedata
	wire         mm_interconnect_0_oct_s1_chipselect;                        // mm_interconnect_0:oct_s1_chipselect -> oct:chipselect
	wire  [31:0] mm_interconnect_0_oct_s1_readdata;                          // oct:readdata -> mm_interconnect_0:oct_s1_readdata
	wire   [1:0] mm_interconnect_0_oct_s1_address;                           // mm_interconnect_0:oct_s1_address -> oct:address
	wire         mm_interconnect_0_oct_s1_write;                             // mm_interconnect_0:oct_s1_write -> oct:write_n
	wire  [31:0] mm_interconnect_0_oct_s1_writedata;                         // mm_interconnect_0:oct_s1_writedata -> oct:writedata
	wire         mm_interconnect_0_waveform_s1_chipselect;                   // mm_interconnect_0:waveform_s1_chipselect -> waveform:chipselect
	wire  [31:0] mm_interconnect_0_waveform_s1_readdata;                     // waveform:readdata -> mm_interconnect_0:waveform_s1_readdata
	wire   [1:0] mm_interconnect_0_waveform_s1_address;                      // mm_interconnect_0:waveform_s1_address -> waveform:address
	wire         mm_interconnect_0_waveform_s1_write;                        // mm_interconnect_0:waveform_s1_write -> waveform:write_n
	wire  [31:0] mm_interconnect_0_waveform_s1_writedata;                    // mm_interconnect_0:waveform_s1_writedata -> waveform:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                     // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                      // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;        // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;          // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;           // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;              // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;             // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;         // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                   // i2c_0:intr -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // spi_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [a0:reset_n, a1:reset_n, a2:reset_n, a3:reset_n, amplitude:reset_n, d0:reset_n, d1:reset_n, d2:reset_n, d3:reset_n, hex_digits_pio:reset_n, i2c_0:rst_n, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, keycode1:reset_n, keycode2:reset_n, keycode3:reset_n, keycode:reset_n, leds_pio:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, oct:reset_n, onchip_memory2_0:reset, phase_incr0:reset_n, phase_incr10:reset_n, phase_incr11:reset_n, phase_incr12:reset_n, phase_incr13:reset_n, phase_incr14:reset_n, phase_incr15:reset_n, phase_incr16:reset_n, phase_incr17:reset_n, phase_incr1:reset_n, phase_incr2:reset_n, phase_incr3:reset_n, phase_incr4:reset_n, phase_incr5:reset_n, phase_incr6:reset_n, phase_incr7:reset_n, phase_incr8:reset_n, phase_incr9:reset_n, r0:reset_n, r1:reset_n, r2:reset_n, r3:reset_n, rst_translator:in_reset, s0:reset_n, s1:reset_n, s2:reset_n, s3:reset_n, sdram_pll:reset, spi_0:reset_n, switches:reset_n, sysid_qsys_0:reset_n, timer:reset_n, usb_gpx:reset_n, usb_irq:reset_n, usb_rst:reset_n, waveform:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	finalProject_a0 a0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_a0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_a0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_a0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_a0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_a0_s1_readdata),   //                    .readdata
		.out_port   (a0_external_connection_export)       // external_connection.export
	);

	finalProject_a0 a1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_a1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_a1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_a1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_a1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_a1_s1_readdata),   //                    .readdata
		.out_port   (a1_external_connection_export)       // external_connection.export
	);

	finalProject_a0 a2 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_a2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_a2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_a2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_a2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_a2_s1_readdata),   //                    .readdata
		.out_port   (a2_external_connection_export)       // external_connection.export
	);

	finalProject_a0 a3 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_a3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_a3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_a3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_a3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_a3_s1_readdata),   //                    .readdata
		.out_port   (a3_external_connection_export)       // external_connection.export
	);

	finalProject_amplitude amplitude (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_amplitude_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_amplitude_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_amplitude_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_amplitude_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_amplitude_s1_readdata),   //                    .readdata
		.out_port   (amp_export)                                 // external_connection.export
	);

	finalProject_a0 d0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_d0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_d0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_d0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_d0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_d0_s1_readdata),   //                    .readdata
		.out_port   (d0_external_connection_export)       // external_connection.export
	);

	finalProject_a0 d1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_d1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_d1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_d1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_d1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_d1_s1_readdata),   //                    .readdata
		.out_port   (d1_external_connection_export)       // external_connection.export
	);

	finalProject_a0 d2 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_d2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_d2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_d2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_d2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_d2_s1_readdata),   //                    .readdata
		.out_port   (d2_external_connection_export)       // external_connection.export
	);

	finalProject_a0 d3 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_d3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_d3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_d3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_d3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_d3_s1_readdata),   //                    .readdata
		.out_port   (d3_external_connection_export)       // external_connection.export
	);

	finalProject_amplitude hex_digits_pio (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_hex_digits_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_digits_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_digits_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_digits_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_digits_pio_s1_readdata),   //                    .readdata
		.out_port   (hex_digits_export)                               // external_connection.export
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (16),
		.FIFO_DEPTH_LOG2 (4)
	) i2c_0 (
		.clk       (clk_clk),                               //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset),       //       reset_sink.reset_n
		.intr      (irq_mapper_receiver0_irq),              // interrupt_sender.irq
		.addr      (mm_interconnect_0_i2c_0_csr_address),   //              csr.address
		.read      (mm_interconnect_0_i2c_0_csr_read),      //                 .read
		.write     (mm_interconnect_0_i2c_0_csr_write),     //                 .write
		.writedata (mm_interconnect_0_i2c_0_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_0_i2c_0_csr_readdata),  //                 .readdata
		.sda_in    (i2c_serial_sda_in),                     //       i2c_serial.sda_in
		.scl_in    (i2c_serial_scl_in),                     //                 .scl_in
		.sda_oe    (i2c_serial_sda_oe),                     //                 .sda_oe
		.scl_oe    (i2c_serial_scl_oe),                     //                 .scl_oe
		.src_data  (),                                      //      (terminated)
		.src_valid (),                                      //      (terminated)
		.src_ready (1'b0),                                  //      (terminated)
		.snk_data  (16'b0000000000000000),                  //      (terminated)
		.snk_valid (1'b0),                                  //      (terminated)
		.snk_ready ()                                       //      (terminated)
	);

	finalProject_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	finalProject_key key (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata), //                    .readdata
		.in_port  (key_external_connection_export)     // external_connection.export
	);

	finalProject_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	finalProject_keycode keycode1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_keycode1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode1_s1_readdata),   //                    .readdata
		.out_port   (keycode1_export)                           // external_connection.export
	);

	finalProject_keycode keycode2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_keycode2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode2_s1_readdata),   //                    .readdata
		.out_port   (keycode2_export)                           // external_connection.export
	);

	finalProject_keycode keycode3 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_keycode3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode3_s1_readdata),   //                    .readdata
		.out_port   (keycode3_export)                           // external_connection.export
	);

	finalProject_leds_pio leds_pio (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_leds_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_pio_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                               // external_connection.export
	);

	finalProject_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	finalProject_keycode oct (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_oct_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_oct_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_oct_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_oct_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_oct_s1_readdata),   //                    .readdata
		.out_port   (oct_external_connection_export)       // external_connection.export
	);

	finalProject_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	finalProject_phase_incr0 phase_incr0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr0_s1_readdata),   //                    .readdata
		.out_port   (phase_incr0_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr1_s1_readdata),   //                    .readdata
		.out_port   (phase_incr1_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr10 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr10_s1_readdata),   //                    .readdata
		.out_port   (phase_incr10_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr11 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr11_s1_readdata),   //                    .readdata
		.out_port   (phase_incr11_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr12 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr12_s1_readdata),   //                    .readdata
		.out_port   (phase_incr12_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr13 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr13_s1_readdata),   //                    .readdata
		.out_port   (phase_incr13_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr14 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr14_s1_readdata),   //                    .readdata
		.out_port   (phase_incr14_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr15 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr15_s1_readdata),   //                    .readdata
		.out_port   (phase_incr15_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr16 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr16_s1_readdata),   //                    .readdata
		.out_port   (phase_incr16_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr17 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr17_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr17_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr17_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr17_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr17_s1_readdata),   //                    .readdata
		.out_port   (phase_incr17_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr2_s1_readdata),   //                    .readdata
		.out_port   (phase_incr2_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr3_s1_readdata),   //                    .readdata
		.out_port   (phase_incr3_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr4_s1_readdata),   //                    .readdata
		.out_port   (phase_incr4_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr5_s1_readdata),   //                    .readdata
		.out_port   (phase_incr5_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr6_s1_readdata),   //                    .readdata
		.out_port   (phase_incr6_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr7 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr7_s1_readdata),   //                    .readdata
		.out_port   (phase_incr7_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr8 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr8_s1_readdata),   //                    .readdata
		.out_port   (phase_incr8_external_connection_export)       // external_connection.export
	);

	finalProject_phase_incr0 phase_incr9 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_phase_incr9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_phase_incr9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_phase_incr9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_phase_incr9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_phase_incr9_s1_readdata),   //                    .readdata
		.out_port   (phase_incr9_external_connection_export)       // external_connection.export
	);

	finalProject_a0 r0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r0_s1_readdata),   //                    .readdata
		.out_port   (r0_external_connection_export)       // external_connection.export
	);

	finalProject_a0 r1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r1_s1_readdata),   //                    .readdata
		.out_port   (r1_external_connection_export)       // external_connection.export
	);

	finalProject_a0 r2 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r2_s1_readdata),   //                    .readdata
		.out_port   (r2_external_connection_export)       // external_connection.export
	);

	finalProject_a0 r3 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r3_s1_readdata),   //                    .readdata
		.out_port   (r3_external_connection_export)       // external_connection.export
	);

	finalProject_a0 s0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s0_s1_readdata),   //                    .readdata
		.out_port   (s0_external_connection_export)       // external_connection.export
	);

	finalProject_a0 s1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s1_s1_readdata),   //                    .readdata
		.out_port   (s1_external_connection_export)       // external_connection.export
	);

	finalProject_a0 s2 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s2_s1_readdata),   //                    .readdata
		.out_port   (s2_external_connection_export)       // external_connection.export
	);

	finalProject_a0 s3 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s3_s1_readdata),   //                    .readdata
		.out_port   (s3_external_connection_export)       // external_connection.export
	);

	finalProject_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	finalProject_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk)                                    //                    c1.clk
	);

	finalProject_spi_0 spi_0 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                            //              irq.irq
		.MISO          (spi0_MISO),                                           //         external.export
		.MOSI          (spi0_MOSI),                                           //                 .export
		.SCLK          (spi0_SCLK),                                           //                 .export
		.SS_n          (spi0_SS_n)                                            //                 .export
	);

	finalProject_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	finalProject_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	finalProject_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	finalProject_usb_gpx usb_gpx (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_usb_gpx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_gpx_s1_readdata), //                    .readdata
		.in_port  (usb_gpx_export)                         // external_connection.export
	);

	finalProject_usb_gpx usb_irq (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_usb_irq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_irq_s1_readdata), //                    .readdata
		.in_port  (usb_irq_export)                         // external_connection.export
	);

	finalProject_usb_rst usb_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_usb_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_usb_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_usb_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_usb_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_usb_rst_s1_readdata),   //                    .readdata
		.out_port   (usb_rst_export)                           // external_connection.export
	);

	finalProject_keycode waveform (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_waveform_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_waveform_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_waveform_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_waveform_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_waveform_s1_readdata),   //                    .readdata
		.out_port   (waveform_external_connection_export)       // external_connection.export
	);

	finalProject_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                           //                             sdram_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                         //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.a0_s1_address                                  (mm_interconnect_0_a0_s1_address),                            //                                    a0_s1.address
		.a0_s1_write                                    (mm_interconnect_0_a0_s1_write),                              //                                         .write
		.a0_s1_readdata                                 (mm_interconnect_0_a0_s1_readdata),                           //                                         .readdata
		.a0_s1_writedata                                (mm_interconnect_0_a0_s1_writedata),                          //                                         .writedata
		.a0_s1_chipselect                               (mm_interconnect_0_a0_s1_chipselect),                         //                                         .chipselect
		.a1_s1_address                                  (mm_interconnect_0_a1_s1_address),                            //                                    a1_s1.address
		.a1_s1_write                                    (mm_interconnect_0_a1_s1_write),                              //                                         .write
		.a1_s1_readdata                                 (mm_interconnect_0_a1_s1_readdata),                           //                                         .readdata
		.a1_s1_writedata                                (mm_interconnect_0_a1_s1_writedata),                          //                                         .writedata
		.a1_s1_chipselect                               (mm_interconnect_0_a1_s1_chipselect),                         //                                         .chipselect
		.a2_s1_address                                  (mm_interconnect_0_a2_s1_address),                            //                                    a2_s1.address
		.a2_s1_write                                    (mm_interconnect_0_a2_s1_write),                              //                                         .write
		.a2_s1_readdata                                 (mm_interconnect_0_a2_s1_readdata),                           //                                         .readdata
		.a2_s1_writedata                                (mm_interconnect_0_a2_s1_writedata),                          //                                         .writedata
		.a2_s1_chipselect                               (mm_interconnect_0_a2_s1_chipselect),                         //                                         .chipselect
		.a3_s1_address                                  (mm_interconnect_0_a3_s1_address),                            //                                    a3_s1.address
		.a3_s1_write                                    (mm_interconnect_0_a3_s1_write),                              //                                         .write
		.a3_s1_readdata                                 (mm_interconnect_0_a3_s1_readdata),                           //                                         .readdata
		.a3_s1_writedata                                (mm_interconnect_0_a3_s1_writedata),                          //                                         .writedata
		.a3_s1_chipselect                               (mm_interconnect_0_a3_s1_chipselect),                         //                                         .chipselect
		.amplitude_s1_address                           (mm_interconnect_0_amplitude_s1_address),                     //                             amplitude_s1.address
		.amplitude_s1_write                             (mm_interconnect_0_amplitude_s1_write),                       //                                         .write
		.amplitude_s1_readdata                          (mm_interconnect_0_amplitude_s1_readdata),                    //                                         .readdata
		.amplitude_s1_writedata                         (mm_interconnect_0_amplitude_s1_writedata),                   //                                         .writedata
		.amplitude_s1_chipselect                        (mm_interconnect_0_amplitude_s1_chipselect),                  //                                         .chipselect
		.d0_s1_address                                  (mm_interconnect_0_d0_s1_address),                            //                                    d0_s1.address
		.d0_s1_write                                    (mm_interconnect_0_d0_s1_write),                              //                                         .write
		.d0_s1_readdata                                 (mm_interconnect_0_d0_s1_readdata),                           //                                         .readdata
		.d0_s1_writedata                                (mm_interconnect_0_d0_s1_writedata),                          //                                         .writedata
		.d0_s1_chipselect                               (mm_interconnect_0_d0_s1_chipselect),                         //                                         .chipselect
		.d1_s1_address                                  (mm_interconnect_0_d1_s1_address),                            //                                    d1_s1.address
		.d1_s1_write                                    (mm_interconnect_0_d1_s1_write),                              //                                         .write
		.d1_s1_readdata                                 (mm_interconnect_0_d1_s1_readdata),                           //                                         .readdata
		.d1_s1_writedata                                (mm_interconnect_0_d1_s1_writedata),                          //                                         .writedata
		.d1_s1_chipselect                               (mm_interconnect_0_d1_s1_chipselect),                         //                                         .chipselect
		.d2_s1_address                                  (mm_interconnect_0_d2_s1_address),                            //                                    d2_s1.address
		.d2_s1_write                                    (mm_interconnect_0_d2_s1_write),                              //                                         .write
		.d2_s1_readdata                                 (mm_interconnect_0_d2_s1_readdata),                           //                                         .readdata
		.d2_s1_writedata                                (mm_interconnect_0_d2_s1_writedata),                          //                                         .writedata
		.d2_s1_chipselect                               (mm_interconnect_0_d2_s1_chipselect),                         //                                         .chipselect
		.d3_s1_address                                  (mm_interconnect_0_d3_s1_address),                            //                                    d3_s1.address
		.d3_s1_write                                    (mm_interconnect_0_d3_s1_write),                              //                                         .write
		.d3_s1_readdata                                 (mm_interconnect_0_d3_s1_readdata),                           //                                         .readdata
		.d3_s1_writedata                                (mm_interconnect_0_d3_s1_writedata),                          //                                         .writedata
		.d3_s1_chipselect                               (mm_interconnect_0_d3_s1_chipselect),                         //                                         .chipselect
		.hex_digits_pio_s1_address                      (mm_interconnect_0_hex_digits_pio_s1_address),                //                        hex_digits_pio_s1.address
		.hex_digits_pio_s1_write                        (mm_interconnect_0_hex_digits_pio_s1_write),                  //                                         .write
		.hex_digits_pio_s1_readdata                     (mm_interconnect_0_hex_digits_pio_s1_readdata),               //                                         .readdata
		.hex_digits_pio_s1_writedata                    (mm_interconnect_0_hex_digits_pio_s1_writedata),              //                                         .writedata
		.hex_digits_pio_s1_chipselect                   (mm_interconnect_0_hex_digits_pio_s1_chipselect),             //                                         .chipselect
		.i2c_0_csr_address                              (mm_interconnect_0_i2c_0_csr_address),                        //                                i2c_0_csr.address
		.i2c_0_csr_write                                (mm_interconnect_0_i2c_0_csr_write),                          //                                         .write
		.i2c_0_csr_read                                 (mm_interconnect_0_i2c_0_csr_read),                           //                                         .read
		.i2c_0_csr_readdata                             (mm_interconnect_0_i2c_0_csr_readdata),                       //                                         .readdata
		.i2c_0_csr_writedata                            (mm_interconnect_0_i2c_0_csr_writedata),                      //                                         .writedata
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.key_s1_address                                 (mm_interconnect_0_key_s1_address),                           //                                   key_s1.address
		.key_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                          //                                         .readdata
		.keycode_s1_address                             (mm_interconnect_0_keycode_s1_address),                       //                               keycode_s1.address
		.keycode_s1_write                               (mm_interconnect_0_keycode_s1_write),                         //                                         .write
		.keycode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                      //                                         .readdata
		.keycode_s1_writedata                           (mm_interconnect_0_keycode_s1_writedata),                     //                                         .writedata
		.keycode_s1_chipselect                          (mm_interconnect_0_keycode_s1_chipselect),                    //                                         .chipselect
		.keycode1_s1_address                            (mm_interconnect_0_keycode1_s1_address),                      //                              keycode1_s1.address
		.keycode1_s1_write                              (mm_interconnect_0_keycode1_s1_write),                        //                                         .write
		.keycode1_s1_readdata                           (mm_interconnect_0_keycode1_s1_readdata),                     //                                         .readdata
		.keycode1_s1_writedata                          (mm_interconnect_0_keycode1_s1_writedata),                    //                                         .writedata
		.keycode1_s1_chipselect                         (mm_interconnect_0_keycode1_s1_chipselect),                   //                                         .chipselect
		.keycode2_s1_address                            (mm_interconnect_0_keycode2_s1_address),                      //                              keycode2_s1.address
		.keycode2_s1_write                              (mm_interconnect_0_keycode2_s1_write),                        //                                         .write
		.keycode2_s1_readdata                           (mm_interconnect_0_keycode2_s1_readdata),                     //                                         .readdata
		.keycode2_s1_writedata                          (mm_interconnect_0_keycode2_s1_writedata),                    //                                         .writedata
		.keycode2_s1_chipselect                         (mm_interconnect_0_keycode2_s1_chipselect),                   //                                         .chipselect
		.keycode3_s1_address                            (mm_interconnect_0_keycode3_s1_address),                      //                              keycode3_s1.address
		.keycode3_s1_write                              (mm_interconnect_0_keycode3_s1_write),                        //                                         .write
		.keycode3_s1_readdata                           (mm_interconnect_0_keycode3_s1_readdata),                     //                                         .readdata
		.keycode3_s1_writedata                          (mm_interconnect_0_keycode3_s1_writedata),                    //                                         .writedata
		.keycode3_s1_chipselect                         (mm_interconnect_0_keycode3_s1_chipselect),                   //                                         .chipselect
		.leds_pio_s1_address                            (mm_interconnect_0_leds_pio_s1_address),                      //                              leds_pio_s1.address
		.leds_pio_s1_write                              (mm_interconnect_0_leds_pio_s1_write),                        //                                         .write
		.leds_pio_s1_readdata                           (mm_interconnect_0_leds_pio_s1_readdata),                     //                                         .readdata
		.leds_pio_s1_writedata                          (mm_interconnect_0_leds_pio_s1_writedata),                    //                                         .writedata
		.leds_pio_s1_chipselect                         (mm_interconnect_0_leds_pio_s1_chipselect),                   //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.oct_s1_address                                 (mm_interconnect_0_oct_s1_address),                           //                                   oct_s1.address
		.oct_s1_write                                   (mm_interconnect_0_oct_s1_write),                             //                                         .write
		.oct_s1_readdata                                (mm_interconnect_0_oct_s1_readdata),                          //                                         .readdata
		.oct_s1_writedata                               (mm_interconnect_0_oct_s1_writedata),                         //                                         .writedata
		.oct_s1_chipselect                              (mm_interconnect_0_oct_s1_chipselect),                        //                                         .chipselect
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.phase_incr0_s1_address                         (mm_interconnect_0_phase_incr0_s1_address),                   //                           phase_incr0_s1.address
		.phase_incr0_s1_write                           (mm_interconnect_0_phase_incr0_s1_write),                     //                                         .write
		.phase_incr0_s1_readdata                        (mm_interconnect_0_phase_incr0_s1_readdata),                  //                                         .readdata
		.phase_incr0_s1_writedata                       (mm_interconnect_0_phase_incr0_s1_writedata),                 //                                         .writedata
		.phase_incr0_s1_chipselect                      (mm_interconnect_0_phase_incr0_s1_chipselect),                //                                         .chipselect
		.phase_incr1_s1_address                         (mm_interconnect_0_phase_incr1_s1_address),                   //                           phase_incr1_s1.address
		.phase_incr1_s1_write                           (mm_interconnect_0_phase_incr1_s1_write),                     //                                         .write
		.phase_incr1_s1_readdata                        (mm_interconnect_0_phase_incr1_s1_readdata),                  //                                         .readdata
		.phase_incr1_s1_writedata                       (mm_interconnect_0_phase_incr1_s1_writedata),                 //                                         .writedata
		.phase_incr1_s1_chipselect                      (mm_interconnect_0_phase_incr1_s1_chipselect),                //                                         .chipselect
		.phase_incr10_s1_address                        (mm_interconnect_0_phase_incr10_s1_address),                  //                          phase_incr10_s1.address
		.phase_incr10_s1_write                          (mm_interconnect_0_phase_incr10_s1_write),                    //                                         .write
		.phase_incr10_s1_readdata                       (mm_interconnect_0_phase_incr10_s1_readdata),                 //                                         .readdata
		.phase_incr10_s1_writedata                      (mm_interconnect_0_phase_incr10_s1_writedata),                //                                         .writedata
		.phase_incr10_s1_chipselect                     (mm_interconnect_0_phase_incr10_s1_chipselect),               //                                         .chipselect
		.phase_incr11_s1_address                        (mm_interconnect_0_phase_incr11_s1_address),                  //                          phase_incr11_s1.address
		.phase_incr11_s1_write                          (mm_interconnect_0_phase_incr11_s1_write),                    //                                         .write
		.phase_incr11_s1_readdata                       (mm_interconnect_0_phase_incr11_s1_readdata),                 //                                         .readdata
		.phase_incr11_s1_writedata                      (mm_interconnect_0_phase_incr11_s1_writedata),                //                                         .writedata
		.phase_incr11_s1_chipselect                     (mm_interconnect_0_phase_incr11_s1_chipselect),               //                                         .chipselect
		.phase_incr12_s1_address                        (mm_interconnect_0_phase_incr12_s1_address),                  //                          phase_incr12_s1.address
		.phase_incr12_s1_write                          (mm_interconnect_0_phase_incr12_s1_write),                    //                                         .write
		.phase_incr12_s1_readdata                       (mm_interconnect_0_phase_incr12_s1_readdata),                 //                                         .readdata
		.phase_incr12_s1_writedata                      (mm_interconnect_0_phase_incr12_s1_writedata),                //                                         .writedata
		.phase_incr12_s1_chipselect                     (mm_interconnect_0_phase_incr12_s1_chipselect),               //                                         .chipselect
		.phase_incr13_s1_address                        (mm_interconnect_0_phase_incr13_s1_address),                  //                          phase_incr13_s1.address
		.phase_incr13_s1_write                          (mm_interconnect_0_phase_incr13_s1_write),                    //                                         .write
		.phase_incr13_s1_readdata                       (mm_interconnect_0_phase_incr13_s1_readdata),                 //                                         .readdata
		.phase_incr13_s1_writedata                      (mm_interconnect_0_phase_incr13_s1_writedata),                //                                         .writedata
		.phase_incr13_s1_chipselect                     (mm_interconnect_0_phase_incr13_s1_chipselect),               //                                         .chipselect
		.phase_incr14_s1_address                        (mm_interconnect_0_phase_incr14_s1_address),                  //                          phase_incr14_s1.address
		.phase_incr14_s1_write                          (mm_interconnect_0_phase_incr14_s1_write),                    //                                         .write
		.phase_incr14_s1_readdata                       (mm_interconnect_0_phase_incr14_s1_readdata),                 //                                         .readdata
		.phase_incr14_s1_writedata                      (mm_interconnect_0_phase_incr14_s1_writedata),                //                                         .writedata
		.phase_incr14_s1_chipselect                     (mm_interconnect_0_phase_incr14_s1_chipselect),               //                                         .chipselect
		.phase_incr15_s1_address                        (mm_interconnect_0_phase_incr15_s1_address),                  //                          phase_incr15_s1.address
		.phase_incr15_s1_write                          (mm_interconnect_0_phase_incr15_s1_write),                    //                                         .write
		.phase_incr15_s1_readdata                       (mm_interconnect_0_phase_incr15_s1_readdata),                 //                                         .readdata
		.phase_incr15_s1_writedata                      (mm_interconnect_0_phase_incr15_s1_writedata),                //                                         .writedata
		.phase_incr15_s1_chipselect                     (mm_interconnect_0_phase_incr15_s1_chipselect),               //                                         .chipselect
		.phase_incr16_s1_address                        (mm_interconnect_0_phase_incr16_s1_address),                  //                          phase_incr16_s1.address
		.phase_incr16_s1_write                          (mm_interconnect_0_phase_incr16_s1_write),                    //                                         .write
		.phase_incr16_s1_readdata                       (mm_interconnect_0_phase_incr16_s1_readdata),                 //                                         .readdata
		.phase_incr16_s1_writedata                      (mm_interconnect_0_phase_incr16_s1_writedata),                //                                         .writedata
		.phase_incr16_s1_chipselect                     (mm_interconnect_0_phase_incr16_s1_chipselect),               //                                         .chipselect
		.phase_incr17_s1_address                        (mm_interconnect_0_phase_incr17_s1_address),                  //                          phase_incr17_s1.address
		.phase_incr17_s1_write                          (mm_interconnect_0_phase_incr17_s1_write),                    //                                         .write
		.phase_incr17_s1_readdata                       (mm_interconnect_0_phase_incr17_s1_readdata),                 //                                         .readdata
		.phase_incr17_s1_writedata                      (mm_interconnect_0_phase_incr17_s1_writedata),                //                                         .writedata
		.phase_incr17_s1_chipselect                     (mm_interconnect_0_phase_incr17_s1_chipselect),               //                                         .chipselect
		.phase_incr2_s1_address                         (mm_interconnect_0_phase_incr2_s1_address),                   //                           phase_incr2_s1.address
		.phase_incr2_s1_write                           (mm_interconnect_0_phase_incr2_s1_write),                     //                                         .write
		.phase_incr2_s1_readdata                        (mm_interconnect_0_phase_incr2_s1_readdata),                  //                                         .readdata
		.phase_incr2_s1_writedata                       (mm_interconnect_0_phase_incr2_s1_writedata),                 //                                         .writedata
		.phase_incr2_s1_chipselect                      (mm_interconnect_0_phase_incr2_s1_chipselect),                //                                         .chipselect
		.phase_incr3_s1_address                         (mm_interconnect_0_phase_incr3_s1_address),                   //                           phase_incr3_s1.address
		.phase_incr3_s1_write                           (mm_interconnect_0_phase_incr3_s1_write),                     //                                         .write
		.phase_incr3_s1_readdata                        (mm_interconnect_0_phase_incr3_s1_readdata),                  //                                         .readdata
		.phase_incr3_s1_writedata                       (mm_interconnect_0_phase_incr3_s1_writedata),                 //                                         .writedata
		.phase_incr3_s1_chipselect                      (mm_interconnect_0_phase_incr3_s1_chipselect),                //                                         .chipselect
		.phase_incr4_s1_address                         (mm_interconnect_0_phase_incr4_s1_address),                   //                           phase_incr4_s1.address
		.phase_incr4_s1_write                           (mm_interconnect_0_phase_incr4_s1_write),                     //                                         .write
		.phase_incr4_s1_readdata                        (mm_interconnect_0_phase_incr4_s1_readdata),                  //                                         .readdata
		.phase_incr4_s1_writedata                       (mm_interconnect_0_phase_incr4_s1_writedata),                 //                                         .writedata
		.phase_incr4_s1_chipselect                      (mm_interconnect_0_phase_incr4_s1_chipselect),                //                                         .chipselect
		.phase_incr5_s1_address                         (mm_interconnect_0_phase_incr5_s1_address),                   //                           phase_incr5_s1.address
		.phase_incr5_s1_write                           (mm_interconnect_0_phase_incr5_s1_write),                     //                                         .write
		.phase_incr5_s1_readdata                        (mm_interconnect_0_phase_incr5_s1_readdata),                  //                                         .readdata
		.phase_incr5_s1_writedata                       (mm_interconnect_0_phase_incr5_s1_writedata),                 //                                         .writedata
		.phase_incr5_s1_chipselect                      (mm_interconnect_0_phase_incr5_s1_chipselect),                //                                         .chipselect
		.phase_incr6_s1_address                         (mm_interconnect_0_phase_incr6_s1_address),                   //                           phase_incr6_s1.address
		.phase_incr6_s1_write                           (mm_interconnect_0_phase_incr6_s1_write),                     //                                         .write
		.phase_incr6_s1_readdata                        (mm_interconnect_0_phase_incr6_s1_readdata),                  //                                         .readdata
		.phase_incr6_s1_writedata                       (mm_interconnect_0_phase_incr6_s1_writedata),                 //                                         .writedata
		.phase_incr6_s1_chipselect                      (mm_interconnect_0_phase_incr6_s1_chipselect),                //                                         .chipselect
		.phase_incr7_s1_address                         (mm_interconnect_0_phase_incr7_s1_address),                   //                           phase_incr7_s1.address
		.phase_incr7_s1_write                           (mm_interconnect_0_phase_incr7_s1_write),                     //                                         .write
		.phase_incr7_s1_readdata                        (mm_interconnect_0_phase_incr7_s1_readdata),                  //                                         .readdata
		.phase_incr7_s1_writedata                       (mm_interconnect_0_phase_incr7_s1_writedata),                 //                                         .writedata
		.phase_incr7_s1_chipselect                      (mm_interconnect_0_phase_incr7_s1_chipselect),                //                                         .chipselect
		.phase_incr8_s1_address                         (mm_interconnect_0_phase_incr8_s1_address),                   //                           phase_incr8_s1.address
		.phase_incr8_s1_write                           (mm_interconnect_0_phase_incr8_s1_write),                     //                                         .write
		.phase_incr8_s1_readdata                        (mm_interconnect_0_phase_incr8_s1_readdata),                  //                                         .readdata
		.phase_incr8_s1_writedata                       (mm_interconnect_0_phase_incr8_s1_writedata),                 //                                         .writedata
		.phase_incr8_s1_chipselect                      (mm_interconnect_0_phase_incr8_s1_chipselect),                //                                         .chipselect
		.phase_incr9_s1_address                         (mm_interconnect_0_phase_incr9_s1_address),                   //                           phase_incr9_s1.address
		.phase_incr9_s1_write                           (mm_interconnect_0_phase_incr9_s1_write),                     //                                         .write
		.phase_incr9_s1_readdata                        (mm_interconnect_0_phase_incr9_s1_readdata),                  //                                         .readdata
		.phase_incr9_s1_writedata                       (mm_interconnect_0_phase_incr9_s1_writedata),                 //                                         .writedata
		.phase_incr9_s1_chipselect                      (mm_interconnect_0_phase_incr9_s1_chipselect),                //                                         .chipselect
		.r0_s1_address                                  (mm_interconnect_0_r0_s1_address),                            //                                    r0_s1.address
		.r0_s1_write                                    (mm_interconnect_0_r0_s1_write),                              //                                         .write
		.r0_s1_readdata                                 (mm_interconnect_0_r0_s1_readdata),                           //                                         .readdata
		.r0_s1_writedata                                (mm_interconnect_0_r0_s1_writedata),                          //                                         .writedata
		.r0_s1_chipselect                               (mm_interconnect_0_r0_s1_chipselect),                         //                                         .chipselect
		.r1_s1_address                                  (mm_interconnect_0_r1_s1_address),                            //                                    r1_s1.address
		.r1_s1_write                                    (mm_interconnect_0_r1_s1_write),                              //                                         .write
		.r1_s1_readdata                                 (mm_interconnect_0_r1_s1_readdata),                           //                                         .readdata
		.r1_s1_writedata                                (mm_interconnect_0_r1_s1_writedata),                          //                                         .writedata
		.r1_s1_chipselect                               (mm_interconnect_0_r1_s1_chipselect),                         //                                         .chipselect
		.r2_s1_address                                  (mm_interconnect_0_r2_s1_address),                            //                                    r2_s1.address
		.r2_s1_write                                    (mm_interconnect_0_r2_s1_write),                              //                                         .write
		.r2_s1_readdata                                 (mm_interconnect_0_r2_s1_readdata),                           //                                         .readdata
		.r2_s1_writedata                                (mm_interconnect_0_r2_s1_writedata),                          //                                         .writedata
		.r2_s1_chipselect                               (mm_interconnect_0_r2_s1_chipselect),                         //                                         .chipselect
		.r3_s1_address                                  (mm_interconnect_0_r3_s1_address),                            //                                    r3_s1.address
		.r3_s1_write                                    (mm_interconnect_0_r3_s1_write),                              //                                         .write
		.r3_s1_readdata                                 (mm_interconnect_0_r3_s1_readdata),                           //                                         .readdata
		.r3_s1_writedata                                (mm_interconnect_0_r3_s1_writedata),                          //                                         .writedata
		.r3_s1_chipselect                               (mm_interconnect_0_r3_s1_chipselect),                         //                                         .chipselect
		.s0_s1_address                                  (mm_interconnect_0_s0_s1_address),                            //                                    s0_s1.address
		.s0_s1_write                                    (mm_interconnect_0_s0_s1_write),                              //                                         .write
		.s0_s1_readdata                                 (mm_interconnect_0_s0_s1_readdata),                           //                                         .readdata
		.s0_s1_writedata                                (mm_interconnect_0_s0_s1_writedata),                          //                                         .writedata
		.s0_s1_chipselect                               (mm_interconnect_0_s0_s1_chipselect),                         //                                         .chipselect
		.s1_s1_address                                  (mm_interconnect_0_s1_s1_address),                            //                                    s1_s1.address
		.s1_s1_write                                    (mm_interconnect_0_s1_s1_write),                              //                                         .write
		.s1_s1_readdata                                 (mm_interconnect_0_s1_s1_readdata),                           //                                         .readdata
		.s1_s1_writedata                                (mm_interconnect_0_s1_s1_writedata),                          //                                         .writedata
		.s1_s1_chipselect                               (mm_interconnect_0_s1_s1_chipselect),                         //                                         .chipselect
		.s2_s1_address                                  (mm_interconnect_0_s2_s1_address),                            //                                    s2_s1.address
		.s2_s1_write                                    (mm_interconnect_0_s2_s1_write),                              //                                         .write
		.s2_s1_readdata                                 (mm_interconnect_0_s2_s1_readdata),                           //                                         .readdata
		.s2_s1_writedata                                (mm_interconnect_0_s2_s1_writedata),                          //                                         .writedata
		.s2_s1_chipselect                               (mm_interconnect_0_s2_s1_chipselect),                         //                                         .chipselect
		.s3_s1_address                                  (mm_interconnect_0_s3_s1_address),                            //                                    s3_s1.address
		.s3_s1_write                                    (mm_interconnect_0_s3_s1_write),                              //                                         .write
		.s3_s1_readdata                                 (mm_interconnect_0_s3_s1_readdata),                           //                                         .readdata
		.s3_s1_writedata                                (mm_interconnect_0_s3_s1_writedata),                          //                                         .writedata
		.s3_s1_chipselect                               (mm_interconnect_0_s3_s1_chipselect),                         //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                         //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                           //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                            //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                        //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                       //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                      //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                     //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                      //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),              //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                 //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),             //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),            //                                         .writedata
		.spi_0_spi_control_port_address                 (mm_interconnect_0_spi_0_spi_control_port_address),           //                   spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                   (mm_interconnect_0_spi_0_spi_control_port_write),             //                                         .write
		.spi_0_spi_control_port_read                    (mm_interconnect_0_spi_0_spi_control_port_read),              //                                         .read
		.spi_0_spi_control_port_readdata                (mm_interconnect_0_spi_0_spi_control_port_readdata),          //                                         .readdata
		.spi_0_spi_control_port_writedata               (mm_interconnect_0_spi_0_spi_control_port_writedata),         //                                         .writedata
		.spi_0_spi_control_port_chipselect              (mm_interconnect_0_spi_0_spi_control_port_chipselect),        //                                         .chipselect
		.switches_s1_address                            (mm_interconnect_0_switches_s1_address),                      //                              switches_s1.address
		.switches_s1_readdata                           (mm_interconnect_0_switches_s1_readdata),                     //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),       //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),      //                                         .readdata
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                         //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                           //                                         .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                        //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                       //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect),                      //                                         .chipselect
		.usb_gpx_s1_address                             (mm_interconnect_0_usb_gpx_s1_address),                       //                               usb_gpx_s1.address
		.usb_gpx_s1_readdata                            (mm_interconnect_0_usb_gpx_s1_readdata),                      //                                         .readdata
		.usb_irq_s1_address                             (mm_interconnect_0_usb_irq_s1_address),                       //                               usb_irq_s1.address
		.usb_irq_s1_readdata                            (mm_interconnect_0_usb_irq_s1_readdata),                      //                                         .readdata
		.usb_rst_s1_address                             (mm_interconnect_0_usb_rst_s1_address),                       //                               usb_rst_s1.address
		.usb_rst_s1_write                               (mm_interconnect_0_usb_rst_s1_write),                         //                                         .write
		.usb_rst_s1_readdata                            (mm_interconnect_0_usb_rst_s1_readdata),                      //                                         .readdata
		.usb_rst_s1_writedata                           (mm_interconnect_0_usb_rst_s1_writedata),                     //                                         .writedata
		.usb_rst_s1_chipselect                          (mm_interconnect_0_usb_rst_s1_chipselect),                    //                                         .chipselect
		.waveform_s1_address                            (mm_interconnect_0_waveform_s1_address),                      //                              waveform_s1.address
		.waveform_s1_write                              (mm_interconnect_0_waveform_s1_write),                        //                                         .write
		.waveform_s1_readdata                           (mm_interconnect_0_waveform_s1_readdata),                     //                                         .readdata
		.waveform_s1_writedata                          (mm_interconnect_0_waveform_s1_writedata),                    //                                         .writedata
		.waveform_s1_chipselect                         (mm_interconnect_0_waveform_s1_chipselect)                    //                                         .chipselect
	);

	finalProject_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
