// finalProject_subsystemA_0.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module finalProject_subsystemA_0 (
	);

endmodule
